

module ula(In1, In2, OP, result, Zero_flag);
	input wire [31:0] In1, In2;
	input wire [3:0] OP;
	output wire [31:0] result;
	output wire Zero_flag;

endmodule
